
module RISCV_Branch_Predictor (
    input brachSignal,
    output brachAddress
);


    
endmodule